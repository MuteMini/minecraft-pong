library ieee;
use ieee.std_logic_1164.all;

ENTITY Registers_tb IS
END Registers_tb;

ARCHITECTURE behaviour IS
    --component
END behaviour;